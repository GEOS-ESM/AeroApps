netcdf sample1 {
dimensions:
	nbatches = UNLIMITED ; // (1 currently)
	batchlen = 1000 ;
	nkt = 7 ;
	nkx = 87 ;
	nqcx = 100 ;
	ndays = 255 ;
	nsyn = 4 ;
	strlen = 50 ;

variables:
	char kt_names(nkt, strlen) ;
		kt_names:name = "Name of GEOS/DAS data types" ;
	char kt_units(nkt, strlen) ;
		kt_units:name = "Units for each GEOS/DAS data type" ;
	char kx_names(nkx, strlen) ;
		kx_names:name = "Name of GEOS/DAS data sources" ;
	char kx_meta(nkx, strlen) ;
		kx_meta:name = "kx specific metadata information" ;
	char qcx_names(nqcx, strlen) ;
		qcx_names:name = "Meaning of each possible value of the quality control exclusion mark" ;
	short lat(nbatches, batchlen) ;
		lat:name = "Latitude" ;
		lat:units = "degrees north" ;
		lat:valid_range = -90.f, 90.f ;
		lat:scale_factor = 0.0099999998f ;
	short lon(nbatches, batchlen) ;
		lon:name = "Longitude" ;
		lon:units = "degrees east" ;
		lon:value_at_90E = 90.f ;
		lon:value_at_90W = -90.f ;
		lon:valid_range = -180.f, 180.f ;
		lon:scale_factor = 0.0099999998f ;
	float lev(nbatches, batchlen) ;
		lev:name = "Pressure level or channel" ;
		lev:units = "hPa or none" ;
	short time(nbatches, batchlen) ;
		time:name = "minutes since 0:00 GMT of first julian day on file" ;
		time:units = "minutes since 1968-05-23 00:00:00.0" ;
		time:add_offset = 32587 ;
		time:valid_range = -180, 65354 ;
	byte kt(nbatches, batchlen) ;
		kt:name = "Data type index" ;
		kt:add_offset = 1 ;
		kt:valid_range = 1, 7 ;
	short kx(nbatches, batchlen) ;
		kx:name = "Data source index" ;
		kx:add_offset = 32768 ;
		kx:valid_range = 1, 87 ;
	long ks(nbatches, batchlen) ;
		ks:name = "Sounding index" ;
		ks:add_offset = 0 ;
		ks:valid_range = 1, 1073741824 ;
	float xm(nbatches, batchlen) ;
		xm:name = "Metadata" ;
		xm:missing_value = 9.9999999e+14f ;
	float obs(nbatches, batchlen) ;
		obs:name = "Observation value" ;
		obs:missing_value = 9.9999999e+14f ;
	byte qcexcl(nbatches, batchlen) ;
		qcexcl:name = "Quality control exclusion mark" ;
		qcexcl:valid_range = 0, 255 ;
	short qchist(nbatches, batchlen) ;
		qchist:name = "Quality control history mark" ;
		qchist:add_offset = 32767 ;
		qchist:valid_range = 0, 65534 ;
	long days(ndays) ;
	long syn_beg(ndays, nsyn) ;
		syn_beg:name = "Begining of synoptic hour for each day" ;
		syn_beg:reference_date = "1968-05-23" ;
		syn_beg:value_at_reference_date = 2440000 ;
		syn_beg:first_julian_day = 2440000 ;
		syn_beg:latest_julian_day = 2440005 ;
		syn_beg:latest_synoptic_hour = 18 ;
	long syn_len(ndays, nsyn) ;
		syn_len:name = "Number of observations for syn. time" ;

// global attributes:
		:source = "Data Assimilation Office, Code 910.3, NASA/GSFC" ;
		:title = "GEOS DAS Observational Data Stream (ODS) File" ;
		:type = "pre_analysis" ;
		:version = "2.02" ;
		:data_info = "Contact data@dao.gsfc.nasa.gov" ;
		:history = "test1                                                                                                                                                                               " ;

data:

 kt_names =
  "surface pressure $                                ",
  "surface u-wind component $                        ",
  "surface v-wind component $                        ",
  "geopotential height $                             ",
  "humidity (dew point) $                            ",
  "u-wind component $                                ",
  "v-wind component $                                " ;

 kt_units =
  "HPa $                                             ",
  "m/s $                                             ",
  "m/s $                                             ",
  "m $                                               ",
  "K $                                               ",
  "m/s $                                             ",
  "m/s $                                             " ;

 kx_names =
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "rawindsonde $                                     ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "tovC $                                            " ;

 kx_meta =
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "oms_file:rawind.oms $                             ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "oms_file:tovC.oms $                               " ;

 qcx_names =
  "valid $                                           ",
  "warning $                                         ",
  "rejected by gross check $                         ",
  "rejected by buddy check $                         ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  " ;

 lat =
  3012, 0, 0, 3012, 0, 3012, 3012, 0, 0, 4582, 0, 0, 0, 0, 4582, 4582, 4582, 
    0, 0, 4582, 3012, 3012, 3012, 3012, 0, 3012, 3012, 0, 0, 4582, 0, 0, 
    4582, 0, 4582, 4582, 4582, 0, 0, 4582, 1051, 0, 1051, 0, 1051, 3012, 
    3012, 3012, 3012, 0, 3012, 3012, 0, 0, 4582, 0, 0, 4582, 0, 4582, 4582, 
    4582, 0, 0, 4582, 1051, 0, 1051, 0, 1051, 3012, 0, 0, 3012, 0, 3012, 
    3012, 0, 0, 4582, 0, 0, 0, 0, 4582, 4582, 4582, 0, 0, 4582, 3012, 3012, 
    3012, 3012, 0, 3012, 3012, 0, 0, 4582, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767 ;

 lon =
  -8090, 0, 0, -8090, 0, -8090, -8090, 0, 0, 10090, 0, 0, 0, 0, 10090, 10090, 
    10090, 0, 0, 10090, -8090, -8090, -8090, -8090, 0, -8090, -8090, 0, 0, 
    10090, 0, 0, 10090, 0, 10090, 10090, 10090, 0, 0, 10090, -7144, 0, -7044, 
    0, -7044, -8090, -8090, -8090, -8090, 0, -8090, -8090, 0, 0, 10090, 0, 0, 
    10090, 0, 10090, 10090, 10090, 0, 0, 10090, -7144, 0, -7044, 0, -7044, 
    -8090, 0, 0, -8090, 0, -8090, -8090, 0, 0, 10090, 0, 0, 0, 0, 10090, 
    10090, 10090, 0, 0, 10090, -8090, -8090, -8090, -8090, 0, -8090, -8090, 
    0, 0, 10090, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767 ;

 lev =
  500 , 0 , 0 , 300 , 0 , 300 , 300 , 0 , 0 , 850 , 0 , 0 , 0 , 0 , 500 , 
    500 , 500 , 0 , 0 , 300 , 500 , 500 , 500 , 300 , 0 , 300 , 300 , 0 , 0 , 
    850 , 0 , 0 , 850 , 0 , 500 , 500 , 500 , 0 , 0 , 300 , 850 , 0 , 700 , 
    0 , 500 , 500 , 500 , 500 , 300 , 0 , 300 , 300 , 0 , 0 , 850 , 0 , 0 , 
    850 , 0 , 500 , 500 , 500 , 0 , 0 , 300 , 850 , 0 , 700 , 0 , 500 , 500 , 
    0 , 0 , 300 , 0 , 300 , 300 , 0 , 0 , 850 , 0 , 0 , 0 , 0 , 500 , 500 , 
    500 , 0 , 0 , 300 , 500 , 500 , 500 , 300 , 0 , 300 , 300 , 0 , 0 , 850 , 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf ;

 time =
  -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, 
    -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, 
    -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, 
    -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, 
    -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, 
    -31507, -31507, -31507, -31507, -31507, -31507, -31507, -31507, -31507, 
    -31507, -31507, -31507, -31507, -31507, -31507, -31507, -31507, -31507, 
    -31507, -31507, -31507, -31507, -31507, -31507, -31507, -32587, -32587, 
    -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, 
    -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, -32587, 
    -24307, -24307, -24307, -24307, -24307, -24307, -24307, -24307, -24307, 
    -24307, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767 ;

 kt =
  3, 0, 0, 3, 0, 4, 4, 0, 0, 3, 0, 0, 0, 0, 5, 6, 4, 0, 0, 3, 3, 4, 5, 3, 0, 
    4, 5, 0, 0, 3, 0, 0, 4, 0, 5, 6, 4, 0, 0, 3, 3, 0, 3, 0, 3, 3, 4, 5, 3, 
    0, 4, 5, 0, 0, 3, 0, 0, 4, 0, 5, 6, 4, 0, 0, 3, 3, 0, 3, 0, 3, 3, 0, 0, 
    3, 0, 4, 4, 0, 0, 3, 0, 0, 0, 0, 5, 6, 4, 0, 0, 3, 3, 4, 5, 3, 0, 4, 5, 
    0, 0, 3, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129 ;

 kx =
  -32761, -32767, -32767, -32761, -32767, -32761, -32761, -32767, -32767, 
    -32761, -32767, -32767, -32767, -32767, -32761, -32761, -32761, -32767, 
    -32767, -32761, -32761, -32761, -32761, -32761, -32767, -32761, -32761, 
    -32767, -32767, -32761, -32767, -32767, -32761, -32767, -32761, -32761, 
    -32761, -32767, -32767, -32761, -32761, -32767, -32761, -32767, -32761, 
    -32761, -32761, -32761, -32761, -32767, -32761, -32761, -32767, -32767, 
    -32761, -32767, -32767, -32761, -32767, -32761, -32761, -32761, -32767, 
    -32767, -32761, -32761, -32767, -32761, -32767, -32761, -32761, -32767, 
    -32767, -32761, -32767, -32761, -32761, -32767, -32767, -32761, -32767, 
    -32767, -32767, -32767, -32761, -32761, -32761, -32767, -32767, -32761, 
    -32761, -32761, -32761, -32761, -32767, -32761, -32761, -32767, -32767, 
    -32761, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767 ;

 xm =
  1.1 , 0 , 0 , 2.2 , 0 , 5 , 22.01 , 0 , 0 , -2.1 , 0 , 0 , 0 , 0 , 33 , 
    21 , 1.05 , 0 , 0 , 0.1 , 2.01 , 1.2 , 4 , 7.1 , 0 , 15.1 , 21.01 , 0 , 
    0 , 14 , 0 , 0 , 66.02 , 0 , 6.2 , 1.1 , 13.7 , 0 , 0 , 1 , 4 , 0 , 
    -6.21 , 0 , 5.11 , 2.01 , 1.2 , 4 , 7.1 , 0 , 15.1 , 21.01 , 0 , 0 , 14 , 
    0 , 0 , 66.02 , 0 , 6.2 , 1.1 , 13.7 , 0 , 0 , 1 , 4 , 0 , -6.21 , 0 , 
    5.11 , 1.1 , 0 , 0 , 2.2 , 0 , 5 , 22.01 , 0 , 0 , -2.1 , 0 , 0 , 0 , 0 , 
    33 , 21 , 1.05 , 0 , 0 , 0.1 , 1.5 , 2.5 , 3.5 , 4.5 , 0 , 6.5 , 7.5 , 
    0 , 0 , 10.5 , FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf ;

 obs =
  5432 , 0 , 0 , 9522 , 0 , 22 , 15 , 0 , 0 , 1524 , 0 , 0 , 0 , 0 , 17 , 
    13 , 268 , 0 , 0 , 9522 , 5371 , 12 , 18 , 9485 , 0 , 28 , 6 , 0 , 0 , 
    1492 , 0 , 0 , 281 , 0 , 21 , 18 , 274 , 0 , 0 , 9355 , 1655 , 0 , 2985 , 
    0 , 5850 , 5371 , 12 , 18 , 9485 , 0 , 28 , 6 , 0 , 0 , 1492 , 0 , 0 , 
    281 , 0 , 21 , 18 , 274 , 0 , 0 , 9355 , 1655 , 0 , 2985 , 0 , 5850 , 
    5432 , 0 , 0 , 9522 , 0 , 22 , 15 , 0 , 0 , 1524 , 0 , 0 , 0 , 0 , 17 , 
    13 , 268 , 0 , 0 , 9522 , 5263 , 15 , 11 , 9376 , 0 , 17 , 22 , 0 , 0 , 
    1367 , FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf ;

 qcexcl =
  2, 0, 0, 3, 0, 1, 4, 0, 0, 1, 0, 0, 0, 0, 2, 1, 4, 0, 0, 1, 0, 1, 0, 1, 0, 
    2, 0, 0, 0, 1, 0, 0, 1, 0, 1, 3, 1, 0, 0, 2, 1, 0, 4, 0, 1, 0, 1, 0, 1, 
    0, 2, 0, 0, 0, 1, 0, 0, 1, 0, 1, 3, 1, 0, 0, 2, 1, 0, 4, 0, 1, 2, 0, 0, 
    3, 0, 1, 4, 0, 0, 1, 0, 0, 0, 0, 2, 1, 4, 0, 0, 1, 1, 2, 2, 5, 0, 7, 2, 
    0, 0, 0, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129 ;

 qchist =
  -32762, -32767, -32767, -32765, -32767, -32750, -32766, -32767, -32767, 
    -32567, -32767, -32767, -32767, -32767, -32751, -32763, -32765, -32767, 
    -32767, -32759, -32765, -32760, -32765, -32744, -32767, -32765, -32760, 
    -32767, -32767, -32765, -32767, -32767, -32752, -32767, -32745, -32749, 
    -32692, -32767, -32767, -32752, -32748, -32767, -32745, -32767, -32723, 
    -32765, -32760, -32765, -32744, -32767, -32765, -32760, -32767, -32767, 
    -32765, -32767, -32767, -32752, -32767, -32745, -32749, -32692, -32767, 
    -32767, -32752, -32748, -32767, -32745, -32767, -32723, -32762, -32767, 
    -32767, -32765, -32767, -32750, -32766, -32767, -32767, -32567, -32767, 
    -32767, -32767, -32767, -32751, -32763, -32765, -32767, -32767, -32759, 
    -32756, -32745, -32734, -32723, -32767, -32701, -32690, -32767, -32767, 
    -32656, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767 ;

 days = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 syn_beg =
  1, 46, 46, 46,
  91, 91, 91, 91,
  91, 91, 91, 91,
  91, 91, 91, 91,
  91, 91, 91, 91,
  91, 91, 91, 91,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101 ;

 syn_len =
  45, 0, 0, 45,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 10,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0 ;
}
