netcdf sample2 {
dimensions:
	nbatches = UNLIMITED ; // (1 currently)
	batchlen = 1000 ;
	ktmax = 7 ;
	kxmax = 87 ;
	ndays = 255 ;
	nsyn = 4 ;
	strlen = 50 ;

variables:
	char kt_names(ktmax, strlen) ;
		kt_names:name = "Name of GEOS/DAS data types" ;
	char kt_units(ktmax, strlen) ;
		kt_units:name = "Units for each GEOS/DAS data type" ;
	char kx_names(kxmax, strlen) ;
		kx_names:name = "Name of GEOS/DAS data sources" ;
	short lat(nbatches, batchlen) ;
		lat:name = "Latitude" ;
		lat:units = "degrees north" ;
		lat:valid_range = -90.f, 90.f ;
		lat:scale_factor = 0.0027466659f ;
	short lon(nbatches, batchlen) ;
		lon:name = "Longitude" ;
		lon:units = "degrees east" ;
		lon:value_at_90E = 90.f ;
		lon:value_at_90W = -90.f ;
		lon:valid_range = -180.f, 180.f ;
		lon:scale_factor = 0.0054933317f ;
	float level(nbatches, batchlen) ;
		level:name = "Pressure level or channel" ;
		level:units = "hPa or none" ;
	short julian(nbatches, batchlen) ;
		julian:name = "Julian day" ;
		julian:reference_date = "1968-05-23$" ;
		julian:value_at_reference_date = 2440000 ;
		julian:add_offset = 17999 ;
		julian:valid_range = 17999, 18254 ;
	short time(nbatches, batchlen) ;
		time:name = "Time stamp since 0 GMT" ;
		time:units = "minutes" ;
		time:valid_range = 0, 1439 ;
	byte kt(nbatches, batchlen) ;
		kt:name = "Data type index" ;
		kt:add_offset = 1 ;
		kt:valid_range = 1, 7 ;
	short kx(nbatches, batchlen) ;
		kx:name = "Data source index" ;
		kx:add_offset = 32768 ;
		kx:valid_range = 1, 87 ;
	short ks(nbatches, batchlen) ;
		ks:name = "Sounding index" ;
		ks:add_offset = 32768 ;
		ks:valid_range = 1, 65535 ;
	long km(nbatches, batchlen) ;
		km:name = "Metadata index" ;
		km:valid_range = 0, 2147483647 ;
		km:missing_value = 0 ;
	float obs(nbatches, batchlen) ;
		obs:name = "Observation value" ;
		obs:missing_value = 9.9999999e+14f ;
	long qc_flag(nbatches, batchlen) ;
		qc_flag:name = "Quality control flag" ;
		qc_flag:add_offset = 32767 ;
		qc_flag:valid_range = 0, 65534 ;
	long days(ndays) ;
	long syn_beg(ndays, nsyn) ;
		syn_beg:name = "Begining of synoptic hour for each day" ;
		syn_beg:reference_date = "1968-05-23$" ;
		syn_beg:value_at_reference_date = 2440000 ;
		syn_beg:first_julian_day = 18000 ;
		syn_beg:latest_julian_day = 18005 ;
		syn_beg:latest_synoptic_hour = 18 ;
	long syn_len(ndays, nsyn) ;
		syn_len:name = "Number of observations for syn. time" ;

// global attributes:
		:source = "Data Assimilation Office, Code 910.3, NASA/GSFC" ;
		:title = "GEOS/DAS Observational Data Stream (ODS) File" ;
		:version = "1.01" ;
		:data_info = "Contact data @dao.gsfc.nasa.gov" ;
		:history = "test1                                                                                                                                                                               " ;

data:

 kt_names =
  "surface pressure $                                ",
  "surface u-wind component $                        ",
  "surface v-wind component $                        ",
  "geopotential height $                             ",
  "humidity (dew point) $                            ",
  "u-wind component $                                ",
  "v-wind component $                                " ;

 kt_units =
  "HPa $                                             ",
  "m/s $                                             ",
  "m/s $                                             ",
  "m $                                               ",
  "K $                                               ",
  "m/s $                                             ",
  "m/s $                                             " ;

 kx_names =
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "rawindsonde $                                     ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "                                                  ",
  "tovC $                                            " ;

 lat =
  10966, 0, 0, 10966, 0, 10966, 10966, 0, 0, 16682, 0, 0, 0, 0, 16682, 16682, 
    16682, 0, 0, 16682, 10966, 10966, 10966, 10966, 0, 10966, 10966, 0, 0, 
    16682, 0, 0, 16682, 0, 16682, 16682, 16682, 0, 0, 16682, 3826, 0, 3826, 
    0, 3826, 10966, 10966, 10966, 10966, 0, 10966, 10966, 0, 0, 16682, 0, 0, 
    16682, 0, 16682, 16682, 16682, 0, 0, 16682, 3826, 0, 3826, 0, 3826, 
    10966, 0, 0, 10966, 0, 10966, 10966, 0, 0, 16682, 0, 0, 0, 0, 16682, 
    16682, 16682, 0, 0, 16682, 10966, 10966, 10966, 10966, 0, 10966, 10966, 
    0, 0, 16682, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767 ;

 lon =
  -14727, 0, 0, -14727, 0, -14727, -14727, 0, 0, 18368, 0, 0, 0, 0, 18368, 
    18368, 18368, 0, 0, 18368, -14727, -14727, -14727, -14727, 0, -14727, 
    -14727, 0, 0, 18368, 0, 0, 18368, 0, 18368, 18368, 18368, 0, 0, 18368, 
    -13005, 0, -12823, 0, -12823, -14727, -14727, -14727, -14727, 0, -14727, 
    -14727, 0, 0, 18368, 0, 0, 18368, 0, 18368, 18368, 18368, 0, 0, 18368, 
    -13005, 0, -12823, 0, -12823, -14727, 0, 0, -14727, 0, -14727, -14727, 0, 
    0, 18368, 0, 0, 0, 0, 18368, 18368, 18368, 0, 0, 18368, -14727, -14727, 
    -14727, -14727, 0, -14727, -14727, 0, 0, 18368, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767 ;

 level =
  500 , 0 , 0 , 300 , 0 , 300 , 300 , 0 , 0 , 850 , 0 , 0 , 0 , 0 , 500 , 
    500 , 500 , 0 , 0 , 300 , 500 , 500 , 500 , 300 , 0 , 300 , 300 , 0 , 0 , 
    850 , 0 , 0 , 850 , 0 , 500 , 500 , 500 , 0 , 0 , 300 , 850 , 0 , 700 , 
    0 , 500 , 500 , 500 , 500 , 300 , 0 , 300 , 300 , 0 , 0 , 850 , 0 , 0 , 
    850 , 0 , 500 , 500 , 500 , 0 , 0 , 300 , 850 , 0 , 700 , 0 , 500 , 500 , 
    0 , 0 , 300 , 0 , 300 , 300 , 0 , 0 , 850 , 0 , 0 , 0 , 0 , 500 , 500 , 
    500 , 0 , 0 , 300 , 500 , 500 , 500 , 300 , 0 , 300 , 300 , 0 , 0 , 850 , 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf ;

 julian =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767 ;

 time =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1080, 1080, 
    1080, 1080, 1080, 1080, 1080, 1080, 1080, 1080, 1080, 1080, 1080, 1080, 
    1080, 1080, 1080, 1080, 1080, 1080, 1080, 1080, 1080, 1080, 1080, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1080, 1080, 1080, 
    1080, 1080, 1080, 1080, 1080, 1080, 1080, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767 ;

 kt =
  3, 0, 0, 3, 0, 4, 4, 0, 0, 3, 0, 0, 0, 0, 5, 6, 4, 0, 0, 3, 3, 4, 5, 3, 0, 
    4, 5, 0, 0, 3, 0, 0, 4, 0, 5, 6, 4, 0, 0, 3, 3, 0, 3, 0, 3, 3, 4, 5, 3, 
    0, 4, 5, 0, 0, 3, 0, 0, 4, 0, 5, 6, 4, 0, 0, 3, 3, 0, 3, 0, 3, 3, 0, 0, 
    3, 0, 4, 4, 0, 0, 3, 0, 0, 0, 0, 5, 6, 4, 0, 0, 3, 3, 4, 5, 3, 0, 4, 5, 
    0, 0, 3, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 
    129, 129, 129, 129, 129 ;

 kx =
  -32761, -32767, -32767, -32761, -32767, -32761, -32761, -32767, -32767, 
    -32761, -32767, -32767, -32767, -32767, -32761, -32761, -32761, -32767, 
    -32767, -32761, -32761, -32761, -32761, -32761, -32767, -32761, -32761, 
    -32767, -32767, -32761, -32767, -32767, -32761, -32767, -32761, -32761, 
    -32761, -32767, -32767, -32761, -32761, -32767, -32761, -32767, -32761, 
    -32761, -32761, -32761, -32761, -32767, -32761, -32761, -32767, -32767, 
    -32761, -32767, -32767, -32761, -32767, -32761, -32761, -32761, -32767, 
    -32767, -32761, -32761, -32767, -32761, -32767, -32761, -32761, -32767, 
    -32767, -32761, -32767, -32761, -32761, -32767, -32767, -32761, -32767, 
    -32767, -32767, -32767, -32761, -32761, -32761, -32767, -32767, -32761, 
    -32761, -32761, -32761, -32761, -32767, -32761, -32761, -32767, -32767, 
    -32761, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, -32767, 
    -32767 ;

 obs =
  5432 , 0 , 0 , 9522 , 0 , 22 , 15 , 0 , 0 , 1524 , 0 , 0 , 0 , 0 , 17 , 
    13 , 268 , 0 , 0 , 9522 , 5371 , 12 , 18 , 9485 , 0 , 28 , 6 , 0 , 0 , 
    1492 , 0 , 0 , 281 , 0 , 21 , 18 , 274 , 0 , 0 , 9355 , 1655 , 0 , 2985 , 
    0 , 5850 , 5371 , 12 , 18 , 9485 , 0 , 28 , 6 , 0 , 0 , 1492 , 0 , 0 , 
    281 , 0 , 21 , 18 , 274 , 0 , 0 , 9355 , 1655 , 0 , 2985 , 0 , 5850 , 
    5432 , 0 , 0 , 9522 , 0 , 22 , 15 , 0 , 0 , 1524 , 0 , 0 , 0 , 0 , 17 , 
    13 , 268 , 0 , 0 , 9522 , 5263 , 15 , 11 , 9376 , 0 , 17 , 22 , 0 , 0 , 
    1367 , FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, FloatInf, 
    FloatInf, FloatInf, FloatInf, FloatInf, FloatInf ;

 qc_flag =
  -32765, -32767, -32767, -32764, -32767, -32766, -32763, -32767, -32767, 
    -32766, -32767, -32767, -32767, -32767, -32765, -32766, -32763, -32767, 
    -32767, -32766, -32767, -32766, -32767, -32766, -32767, -32765, -32767, 
    -32767, -32767, -32766, -32767, -32767, -32766, -32767, -32766, -32764, 
    -32766, -32767, -32767, -32765, -32766, -32767, -32763, -32767, -32766, 
    -32767, -32766, -32767, -32766, -32767, -32765, -32767, -32767, -32767, 
    -32766, -32767, -32767, -32766, -32767, -32766, -32764, -32766, -32767, 
    -32767, -32765, -32766, -32767, -32763, -32767, -32766, -32765, -32767, 
    -32767, -32764, -32767, -32766, -32763, -32767, -32767, -32766, -32767, 
    -32767, -32767, -32767, -32765, -32766, -32763, -32767, -32767, -32766, 
    -32766, -32765, -32765, -32762, -32767, -32760, -32765, -32767, -32767, 
    -32767, -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647, 
    -2147483647, -2147483647, -2147483647, -2147483647, -2147483647 ;

 days = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 syn_beg =
  1, 46, 46, 46,
  91, 91, 91, 91,
  91, 91, 91, 91,
  91, 91, 91, 91,
  91, 91, 91, 91,
  91, 91, 91, 91,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101,
  101, 101, 101, 101 ;

 syn_len =
  45, 0, 0, 45,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 10,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0,
  0, 0, 0, 0 ;
}
